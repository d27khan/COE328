library verilog;
use verilog.vl_types.all;
entity lab1_schm2_vlg_vec_tst is
end lab1_schm2_vlg_vec_tst;
