library verilog;
use verilog.vl_types.all;
entity GPU2_vlg_vec_tst is
end GPU2_vlg_vec_tst;
