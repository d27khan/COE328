library verilog;
use verilog.vl_types.all;
entity LAB2SCHEM2_vlg_vec_tst is
end LAB2SCHEM2_vlg_vec_tst;
