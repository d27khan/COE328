library verilog;
use verilog.vl_types.all;
entity lab1schm_vlg_vec_tst is
end lab1schm_vlg_vec_tst;
