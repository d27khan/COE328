library verilog;
use verilog.vl_types.all;
entity LAB2SCHEM2 is
    port(
        f               : out    vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic
    );
end LAB2SCHEM2;
