library verilog;
use verilog.vl_types.all;
entity Latch2Schem_vlg_vec_tst is
end Latch2Schem_vlg_vec_tst;
