library verilog;
use verilog.vl_types.all;
entity modifiedmux_vlg_vec_tst is
end modifiedmux_vlg_vec_tst;
