library verilog;
use verilog.vl_types.all;
entity Johnsschem_vlg_vec_tst is
end Johnsschem_vlg_vec_tst;
