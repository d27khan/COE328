library verilog;
use verilog.vl_types.all;
entity dec3to8_vlg_check_tst is
    port(
        y0              : in     vl_logic;
        y1              : in     vl_logic;
        y2              : in     vl_logic;
        y3              : in     vl_logic;
        y20             : in     vl_logic;
        y21             : in     vl_logic;
        y22             : in     vl_logic;
        y23             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end dec3to8_vlg_check_tst;
