library verilog;
use verilog.vl_types.all;
entity lab5test_vlg_vec_tst is
end lab5test_vlg_vec_tst;
