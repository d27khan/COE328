library verilog;
use verilog.vl_types.all;
entity Latch1schem_vlg_vec_tst is
end Latch1schem_vlg_vec_tst;
