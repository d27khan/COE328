library verilog;
use verilog.vl_types.all;
entity lab1schm is
    port(
        f               : out    vl_logic;
        x2              : in     vl_logic;
        x3              : in     vl_logic;
        x1              : in     vl_logic
    );
end lab1schm;
