library verilog;
use verilog.vl_types.all;
entity lab1schm_vlg_check_tst is
    port(
        f               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab1schm_vlg_check_tst;
