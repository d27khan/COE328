library verilog;
use verilog.vl_types.all;
entity encode_vlg_vec_tst is
end encode_vlg_vec_tst;
