library verilog;
use verilog.vl_types.all;
entity TEST4to16_vlg_vec_tst is
end TEST4to16_vlg_vec_tst;
