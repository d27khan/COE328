library verilog;
use verilog.vl_types.all;
entity fsmSchem_vlg_vec_tst is
end fsmSchem_vlg_vec_tst;
