library verilog;
use verilog.vl_types.all;
entity MealyFSMschem_vlg_vec_tst is
end MealyFSMschem_vlg_vec_tst;
