library verilog;
use verilog.vl_types.all;
entity test_moore_vlg_vec_tst is
end test_moore_vlg_vec_tst;
