--Author: Daniel Khan (500898010)
--COE318 (Section 041)
--Lab 4:  VHDL for Combinational Circuits and Storage Elements

LIBRARY ieee;								--Defining all libraries and packages
USE ieee.std_logic_1164.all;

ENTITY encod IS 
	PORT( w  : IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- creating a Vector w inputs
			y 	: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);  -- y output vectors
			z  : OUT STD_LOGIC); -- z output
END encod;

ARCHITECTURE Behavior OF encod IS
BEGIN
	PROCESS(w) 
	BEGIN
		y<="00";
		IF w(1) ='1' THEN y<= "01"; END IF; -- encoding all inputs to give a specific output
		IF w(2) ='1' THEN y<= "10"; END IF;
		IF w(3) ='1' THEN y<= "11"; END IF;
		
		z<='1';
		IF w ="0000" THEN z<='0'; END IF;
	END PROCESS;
END Behavior;
