library verilog;
use verilog.vl_types.all;
entity TESTdec3to8_vlg_vec_tst is
end TESTdec3to8_vlg_vec_tst;
