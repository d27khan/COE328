library verilog;
use verilog.vl_types.all;
entity Lab2schm_vlg_vec_tst is
end Lab2schm_vlg_vec_tst;
