library verilog;
use verilog.vl_types.all;
entity ASUa_vlg_vec_tst is
end ASUa_vlg_vec_tst;
