library verilog;
use verilog.vl_types.all;
entity GPU3_vlg_vec_tst is
end GPU3_vlg_vec_tst;
